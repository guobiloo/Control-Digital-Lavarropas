-- Vhdl test bench created from schematic /home/joak/Estudio/electronica digital/tps/TP 2/lavarropas/contadorAs5.sch - Sun Jun 21 20:32:53 2015
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY contadorAs5_contadorAs5_sch_tb IS
END contadorAs5_contadorAs5_sch_tb;
ARCHITECTURE behavioral OF contadorAs5_contadorAs5_sch_tb IS 

   COMPONENT contadorAs5
   PORT( salidaQ	:	OUT	STD_LOGIC; 
          reloj	:	IN	STD_LOGIC);
   END COMPONENT;

   SIGNAL salidaQ	:	STD_LOGIC;
   SIGNAL reloj	:	STD_LOGIC;

BEGIN

   UUT: contadorAs5 PORT MAP(
		salidaQ => salidaQ, 
		reloj => reloj
   );

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
	reloj<='0';
	for it in 0 to 20 loop
		wait for 10 ns;
		reloj<='1';
		wait for 10 ns;
		reloj<='0';
	end loop;
      WAIT; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
